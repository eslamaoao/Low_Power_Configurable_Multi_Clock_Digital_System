module INV
( 
input wire IN,
output wire OUT
);

assign OUT = ~ IN ;
endmodule
